///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SL2_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Input: A (32-bit)
reg[31:0] A;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: S (32-bit)
wire[31:0] S;
///////////////////////////////////////////////////////////////////////////////////

SL2_32 mySE(.I(A), .O(S));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: A=3782
$display("Testing A=3782");
A=3782;   #10; 
verifyEqual32(S, A*4);
////////////////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end

endmodule
